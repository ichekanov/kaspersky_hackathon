component alphabot.Printnum

endpoints {
    printnum : alphabot.Printnum
}